
module pll (
	clk_in_clk,
	clk_out_clk,
	reset_reset);	

	input		clk_in_clk;
	output		clk_out_clk;
	input		reset_reset;
endmodule
